module Comparison(SW, comparisonBinary);

	input SW[9:0];
	
	output comparisonBinary[3:0];
	
	
	
endmodule 
