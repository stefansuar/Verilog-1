module SevenSegment(hexDisplay, HEX0, HEX1);
	input [7:0]hexDisplay;
	output [7:0]HEX0, [7:0]HEX1;
	
	assign hDigit0 = hexDisplay[3:0];
	assign hDigit1 = hexDisplay[7:4];
	
	always @(hexDisplay)
	case (hDigit0)
		4'b0000: HEX0=7'b1111110;
		4'b0001: HEX0=7'b1001111;
		4'b0010: HEX0=7'b0010010;
		4'b0011: HEX0=7'b0000110;
		4'b0100: HEX0=7'b1001100;
		4'b0101: HEX0=7'b0100100;
		4'b0110: HEX0=7'b0100000;
		4'b0111: HEX0=7'b0001111;
		4'b1000: HEX0=7'b0000000;
		4'b1001: HEX0=7'b0000100;
		4'b1010: HEX0=7'b0001000;
		4'b1011: HEX0=7'b1100000;
		4'b1100: HEX0=7'b0110001;
		4'b1101: HEX0=7'b1000010;
		4'b1110: HEX0=7'b0110000;
		4'b1111: HEX0=7'b0111000;
	endcase
	case (hDigit1)
		4'b0000: HEX1=7'b1111110;
		4'b0001: HEX1=7'b1001111;
		4'b0010: HEX1=7'b0010010;
		4'b0011: HEX1=7'b0000110;
		4'b0100: HEX1=7'b1001100;
		4'b0101: HEX1=7'b0100100;
		4'b0110: HEX1=7'b0100000;
		4'b0111: HEX1=7'b0001111;
		4'b1000: HEX1=7'b0000000;
		4'b1001: HEX1=7'b0000100;
		4'b1010: HEX1=7'b0001000;
		4'b1011: HEX1=7'b1100000;
		4'b1100: HEX1=7'b0110001;
		4'b1101: HEX1=7'b1000010;
		4'b1110: HEX1=7'b0110000;
		4'b1111: HEX1=7'b0111000;
	endcase

endmodule 
