module Logical(SW, logicalBinary);

	input SW[9:0];
	
	output logicalBinary[7:0];
	
	
	
endmodule 
