module Arithmetic(SW, arithmeticBinary);

	input SW[9:0];
	
	output arithmeticBinary[8:0];
	
	

endmodule 
